* C:\FOSSEE\eSim\library\SubcircuitLibrary\switch-a\switch-a.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/08/24 16:54:19

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC2  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC2-Pad3_ ? sky130_fd_pr__pfet_01v8		
SC6  Net-_SC5-Pad1_ Net-_SC1-Pad1_ Net-_SC2-Pad3_ ? sky130_fd_pr__pfet_01v8		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ GND ? sky130_fd_pr__nfet_01v8		
SC5  Net-_SC5-Pad1_ Net-_SC1-Pad1_ ? ? sky130_fd_pr__nfet_01v8		
SC4  Net-_SC4-Pad1_ Net-_SC1-Pad1_ ? ? sky130_fd_pr__pfet_01v8		
SC8  Net-_SC3-Pad3_ Net-_SC5-Pad1_ Net-_SC4-Pad1_ ? sky130_fd_pr__pfet_01v8		
SC7  ? Net-_SC5-Pad1_ Net-_SC4-Pad1_ ? sky130_fd_pr__nfet_01v8		
SC3  ? Net-_SC1-Pad1_ Net-_SC3-Pad3_ ? sky130_fd_pr__nfet_01v8		
U1  ? ? ? ? ? PORT		

.end
